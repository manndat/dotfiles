library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_misc.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;

--description of unit (portmap)
entity is
  port (

  );
end;

architecture behavioral of is
--signals

begin
  --processes
  process
  begin

  end process;
end behavioral;
